library verilog;
use verilog.vl_types.all;
entity experiment1_rsp_xbar_mux_001 is
    port(
        sink0_valid     : in     vl_logic;
        sink0_data      : in     vl_logic_vector(89 downto 0);
        sink0_channel   : in     vl_logic_vector(7 downto 0);
        sink0_startofpacket: in     vl_logic;
        sink0_endofpacket: in     vl_logic;
        sink0_ready     : out    vl_logic;
        sink1_valid     : in     vl_logic;
        sink1_data      : in     vl_logic_vector(89 downto 0);
        sink1_channel   : in     vl_logic_vector(7 downto 0);
        sink1_startofpacket: in     vl_logic;
        sink1_endofpacket: in     vl_logic;
        sink1_ready     : out    vl_logic;
        sink2_valid     : in     vl_logic;
        sink2_data      : in     vl_logic_vector(89 downto 0);
        sink2_channel   : in     vl_logic_vector(7 downto 0);
        sink2_startofpacket: in     vl_logic;
        sink2_endofpacket: in     vl_logic;
        sink2_ready     : out    vl_logic;
        sink3_valid     : in     vl_logic;
        sink3_data      : in     vl_logic_vector(89 downto 0);
        sink3_channel   : in     vl_logic_vector(7 downto 0);
        sink3_startofpacket: in     vl_logic;
        sink3_endofpacket: in     vl_logic;
        sink3_ready     : out    vl_logic;
        sink4_valid     : in     vl_logic;
        sink4_data      : in     vl_logic_vector(89 downto 0);
        sink4_channel   : in     vl_logic_vector(7 downto 0);
        sink4_startofpacket: in     vl_logic;
        sink4_endofpacket: in     vl_logic;
        sink4_ready     : out    vl_logic;
        sink5_valid     : in     vl_logic;
        sink5_data      : in     vl_logic_vector(89 downto 0);
        sink5_channel   : in     vl_logic_vector(7 downto 0);
        sink5_startofpacket: in     vl_logic;
        sink5_endofpacket: in     vl_logic;
        sink5_ready     : out    vl_logic;
        sink6_valid     : in     vl_logic;
        sink6_data      : in     vl_logic_vector(89 downto 0);
        sink6_channel   : in     vl_logic_vector(7 downto 0);
        sink6_startofpacket: in     vl_logic;
        sink6_endofpacket: in     vl_logic;
        sink6_ready     : out    vl_logic;
        sink7_valid     : in     vl_logic;
        sink7_data      : in     vl_logic_vector(89 downto 0);
        sink7_channel   : in     vl_logic_vector(7 downto 0);
        sink7_startofpacket: in     vl_logic;
        sink7_endofpacket: in     vl_logic;
        sink7_ready     : out    vl_logic;
        src_valid       : out    vl_logic;
        src_data        : out    vl_logic_vector(89 downto 0);
        src_channel     : out    vl_logic_vector(7 downto 0);
        src_startofpacket: out    vl_logic;
        src_endofpacket : out    vl_logic;
        src_ready       : in     vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
end experiment1_rsp_xbar_mux_001;
